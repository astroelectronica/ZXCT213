.title KiCad schematic
.include "C:/AE/ZXCT213/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/ZXCT213/ZXCT213.LIB"
I1 /IN- 0 DC {ILOAD} 
XU1 /VREF 0 /VSUPPLY /VIN /IN- /CNV ZXCT213
R1 /IN- /VIN {RSNS}
XU2 /OUT 0 CEU4J2X7R2A103K125AE_s
R2 /CNV /OUT {ROUT}
V3 /VSUPPLY 0 DC {VSUPPLY} 
V1 /VIN 0 DC {VIN} 
V2 /VREF 0 DC {VREF} 
.end
